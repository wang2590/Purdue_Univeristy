library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity lab11 is

end;

architecture behavioral of lab11 is
begin

end behavioral;

